<?xml version="1.0" encoding="UTF-8" standalone="yes"?>

<item>
<title>[COLOR yellow]_**_  [/COLOR][COLOR  skyblue] Temporada 1 [/COLOR][COLOR yellow]  _**_[/COLOR]</title>
<link>$doregex[makelist]</link>
<regex>
  <name>makelist</name>
  <listrepeat><![CDATA[
        <title>[COLOR yellow] [makelist.param3] [/COLOR]</title>
        <link>$doregex[getUrl]</link>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
]]></listrepeat>
<expres><![CDATA[href="\/.*,(.*?),list.*\n.*\n.*\n.*href="\/([^"]*)".*?>(.*?)<]]></expres>
<page>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t1-castellano-52961</page>
<cookieJar></cookieJar>
</regex>
<regex>
<name>getUrl</name>
<expres>DownloadUrl":"([^"]+)<expres>
<page>http://diskokosmiko.mx/action/DownloadFile?location=fi&f=[makelist.param1]</page>
<rawpost>fileId=[makelist.param1]&__RequestVerificationToken=$doregex[tok]</rawpost>
<referer>http://diskokosmiko.mx/[makelist.param2]</referer>
<connection>keep-alive</connection>
<accept>*/*</accept>
<X-Req>XMLHttpRequest</X-Req>
<cookieJar></cookieJar>
</regex>
<regex>
<name>tok</name>
<expres>DownloadFile.*RequestVerificationToken.*?value="([^"]+)<expres>
<page>http://diskokosmiko.mx/[makelist.param2]</page>
<referer>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t1-castellano-52961</referer>
<connection>keep-alive</connection>
<cookieJar></cookieJar>
</regex>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
</item>

<item>
<title>[COLOR yellow]_**_  [/COLOR][COLOR  skyblue] Temporada 2 [/COLOR][COLOR yellow]  _**_[/COLOR]</title>
<link>$doregex[makelist]</link>
<regex>
  <name>makelist</name>
  <listrepeat><![CDATA[
        <title>[COLOR yellow] [makelist.param3] [/COLOR]</title>
        <link>$doregex[getUrl]</link>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
]]></listrepeat>
<expres><![CDATA[href="\/.*,(.*?),list.*\n.*\n.*\n.*href="\/([^"]*)".*?>(.*?)<]]></expres>
<page>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t2-castellano-53151</page>
<cookieJar></cookieJar>
</regex>
<regex>
<name>getUrl</name>
<expres>DownloadUrl":"([^"]+)<expres>
<page>http://diskokosmiko.mx/action/DownloadFile?location=fi&f=[makelist.param1]</page>
<rawpost>fileId=[makelist.param1]&__RequestVerificationToken=$doregex[tok]</rawpost>
<referer>http://diskokosmiko.mx/[makelist.param2]</referer>
<connection>keep-alive</connection>
<accept>*/*</accept>
<X-Req>XMLHttpRequest</X-Req>
<cookieJar></cookieJar>
</regex>
<regex>
<name>tok</name>
<expres>DownloadFile.*RequestVerificationToken.*?value="([^"]+)<expres>
<page>http://diskokosmiko.mx/[makelist.param2]</page>
<referer>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t2-castellano-53151</referer>
<connection>keep-alive</connection>
<cookieJar></cookieJar>
</regex>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
</item>

<item>
<title>[COLOR yellow]_**_  [/COLOR][COLOR  skyblue] Temporada 3 [/COLOR][COLOR yellow]  _**_[/COLOR]</title>
<link>$doregex[makelist]</link>
<regex>
  <name>makelist</name>
  <listrepeat><![CDATA[
        <title>[COLOR yellow] [makelist.param3] [/COLOR]</title>
        <link>$doregex[getUrl]</link>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
]]></listrepeat>
<expres><![CDATA[href="\/.*,(.*?),list.*\n.*\n.*\n.*href="\/([^"]*)".*?>(.*?)<]]></expres>
<page>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t3-castellano-53401/list,1,2</page>
<cookieJar></cookieJar>
</regex>
<regex>
<name>getUrl</name>
<expres>DownloadUrl":"([^"]+)<expres>
<page>http://diskokosmiko.mx/action/DownloadFile?location=fi&f=[makelist.param1]</page>
<rawpost>fileId=[makelist.param1]&__RequestVerificationToken=$doregex[tok]</rawpost>
<referer>http://diskokosmiko.mx/[makelist.param2]</referer>
<connection>keep-alive</connection>
<accept>*/*</accept>
<X-Req>XMLHttpRequest</X-Req>
<cookieJar></cookieJar>
</regex>
<regex>
<name>tok</name>
<expres>DownloadFile.*RequestVerificationToken.*?value="([^"]+)<expres>
<page>http://diskokosmiko.mx/[makelist.param2]</page>
<referer>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t3-castellano-53401/list,1,2</referer>
<connection>keep-alive</connection>
<cookieJar></cookieJar>
</regex>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
</item>

<item>
<title>[COLOR yellow]_**_  [/COLOR][COLOR  skyblue] temporada 4 [/COLOR][COLOR yellow]  _**_[/COLOR]</title>
<link>$doregex[makelist]</link>
<regex>
  <name>makelist</name>
  <listrepeat><![CDATA[
        <title>[COLOR yellow] [makelist.param3] [/COLOR]</title>
        <link>$doregex[getUrl]</link>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
]]></listrepeat>
<expres><![CDATA[href="\/.*,(.*?),list.*\n.*\n.*\n.*href="\/([^"]*)".*?>(.*?)<]]></expres>
<page>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t4-castellano-53598</page>
<cookieJar></cookieJar>
</regex>
<regex>
<name>getUrl</name>
<expres>DownloadUrl":"([^"]+)<expres>
<page>http://diskokosmiko.mx/action/DownloadFile?location=fi&f=[makelist.param1]</page>
<rawpost>fileId=[makelist.param1]&__RequestVerificationToken=$doregex[tok]</rawpost>
<referer>http://diskokosmiko.mx/[makelist.param2]</referer>
<connection>keep-alive</connection>
<accept>*/*</accept>
<X-Req>XMLHttpRequest</X-Req>
<cookieJar></cookieJar>
</regex>
<regex>
<name>tok</name>
<expres>DownloadFile.*RequestVerificationToken.*?value="([^"]+)<expres>
<page>http://diskokosmiko.mx/[makelist.param2]</page>
<referer>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t4-castellano-53598</referer>
<connection>keep-alive</connection>
<cookieJar></cookieJar>
</regex>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
</item>

<item>
<title>[COLOR yellow]_**_  [/COLOR][COLOR  skyblue]  [/COLOR][COLOR yellow]  _**_[/COLOR]</title>
<link>$doregex[makelist]</link>
<regex>
  <name>makelist</name>
  <listrepeat><![CDATA[
        <title>[COLOR yellow] [makelist.param3] [/COLOR]</title>
        <link>$doregex[getUrl]</link>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
]]></listrepeat>
<expres><![CDATA[href="\/.*,(.*?),list.*\n.*\n.*\n.*href="\/([^"]*)".*?>(.*?)<]]></expres>
<page></page>
<cookieJar></cookieJar>
</regex>
<regex>
<name>getUrl</name>
<expres>DownloadUrl":"([^"]+)<expres>
<page>http://diskokosmiko.mx/action/DownloadFile?location=fi&f=[makelist.param1]</page>
<rawpost>fileId=[makelist.param1]&__RequestVerificationToken=$doregex[tok]</rawpost>
<referer>http://diskokosmiko.mx/[makelist.param2]</referer>
<connection>keep-alive</connection>
<accept>*/*</accept>
<X-Req>XMLHttpRequest</X-Req>
<cookieJar></cookieJar>
</regex>
<regex>
<name>tok</name>
<expres>DownloadFile.*RequestVerificationToken.*?value="([^"]+)<expres>
<page>http://diskokosmiko.mx/[makelist.param2]</page>
<referer></referer>
<connection>keep-alive</connection>
<cookieJar></cookieJar>
</regex>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
</item>

<item>
<title>[COLOR yellow]_**_  [/COLOR][COLOR  skyblue] Temporada 5 [/COLOR][COLOR yellow]  _**_[/COLOR]</title>
<link>$doregex[makelist]</link>
<regex>
  <name>makelist</name>
  <listrepeat><![CDATA[
        <title>[COLOR yellow] [makelist.param3] [/COLOR]</title>
        <link>$doregex[getUrl]</link>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
]]></listrepeat>
<expres><![CDATA[href="\/.*,(.*?),list.*\n.*\n.*\n.*href="\/([^"]*)".*?>(.*?)<]]></expres>
<page>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t5-castellano-53704</page>
<cookieJar></cookieJar>
</regex>
<regex>
<name>getUrl</name>
<expres>DownloadUrl":"([^"]+)<expres>
<page>http://diskokosmiko.mx/action/DownloadFile?location=fi&f=[makelist.param1]</page>
<rawpost>fileId=[makelist.param1]&__RequestVerificationToken=$doregex[tok]</rawpost>
<referer>http://diskokosmiko.mx/[makelist.param2]</referer>
<connection>keep-alive</connection>
<accept>*/*</accept>
<X-Req>XMLHttpRequest</X-Req>
<cookieJar></cookieJar>
</regex>
<regex>
<name>tok</name>
<expres>DownloadFile.*RequestVerificationToken.*?value="([^"]+)<expres>
<page>http://diskokosmiko.mx/[makelist.param2]</page>
<referer>http://diskokosmiko.mx/gemma-valencia/aqui-no-hay-quien-viva-t5-castellano-53704</referer>
<connection>keep-alive</connection>
<cookieJar></cookieJar>
</regex>
<fanart>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</fanart>
<thumbnail>http://www.seriespapaya.com/uploads/Aqui-no-hay-quien-viva69.jpg</thumbnail>
</item>
